-- VHDL code for stepper drivers
-- Generate clock and watch the safety end stops

-- Autor: Rodolfo Cavour Moretti Schiavi

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_unsigned.all;
use IEEE.NUMERIC_STD.all;

entity stepper_angular is
  port (
    clk_50Mhz : in  std_logic; -- System clock
	 clk_step  : out std_logic :='0'; -- Output clock for the driver generate with this logic
	 velocity_in : in std_logic_vector(3 downto 0) :="0101"; -- velocity_in with 16 options, can be increased
	 distance_in : in integer range 0 to 511 := 50; -- Millimeters that the stepper will move
	 reset : in std_logic := '1' -- Reset for cleaning the variables
	 );
end stepper_angular;

architecture Behavioral of stepper_angular is
	signal state: std_logic :='0'; -- Logic signal for the stepper clock

begin
   PROCESS (clk_50Mhz, velocity_in, reset, distance_in)

   VARIABLE t :INTEGER RANGE 0 TO 2097151:= 0; -- Time counter
	Variable dividend_acel: INTEGER RANGE 0 TO 5000020:= 5000000;	-- Variable to apply aceleration
   CONSTANT dividend :INTEGER RANGE 0 TO 1048575:= 498047;	-- clock divider for 50MHz to reach values within the stepper necessities
	variable distance: integer range 0 to 65535 := distance_in*90; -- Convertion for 1,8 degree stepper and a step 1,75mm/rev
																						-- to change this use the following equation: distance_in*degress*step/360
  

	BEGIN
		IF (clk_50Mhz'EVENT AND clk_50Mhz='1') THEN
			IF (velocity_in > 0) and (distance > 0) and (reset='0') THEN -- Only allows movimentation if the velocity and the distance is greather than 0
				t := t + 1;
				IF (CONV_INTEGER(velocity_in)*t >= dividend_acel) THEN -- This applied logic is used to increase and decrease the clock with the velocity parameter
				   t := 0;
					state <= not state; -- Changes the clk stepper state
					distance := distance - 1; -- Decrease the distance, because on step occured
				END IF;
			END IF;
			IF (dividend_acel > dividend) and (distance > 10) then -- Verify the distance to apply aceleration
					dividend_acel := dividend_acel -1;
			END IF;
			IF(dividend_acel < 5000000) and (distance < 10) then -- Verify the distance to apply the deceleration
				dividend_acel := dividend_acel + 1;
			END IF;
		END IF;
		IF (reset = '1') then -- Reset the distance variable
			distance:=distance_in*90;
		END IF;
	END PROCESS;
	
	-- Apply the signals to the ports
	clk_step<=state;

end Behavioral;