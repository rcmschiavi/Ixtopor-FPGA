-- sopc_2.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sopc_2 is
	port (
		botao_export     : in    std_logic                     := '0';             --     botao.export
		clk_clk          : in    std_logic                     := '0';             --       clk.clk
		entrada_c_export : in    std_logic_vector(7 downto 0)  := (others => '0'); -- entrada_c.export
		hex0_export      : out   std_logic_vector(7 downto 0);                     --      hex0.export
		hex1_export      : out   std_logic_vector(7 downto 0);                     --      hex1.export
		hex2_export      : out   std_logic_vector(7 downto 0);                     --      hex2.export
		hex3_export      : out   std_logic_vector(7 downto 0);                     --      hex3.export
		hex5_export      : out   std_logic_vector(7 downto 0);                     --      hex5.export
		hex_4_export     : out   std_logic_vector(7 downto 0);                     --     hex_4.export
		motor2_export    : out   std_logic_vector(13 downto 0);                    --    motor2.export
		motor3_export    : out   std_logic_vector(13 downto 0);                    --    motor3.export
		motor4_export    : out   std_logic_vector(13 downto 0);                    --    motor4.export
		motor_1_export   : out   std_logic_vector(13 downto 0);                    --   motor_1.export
		porta_a_export   : inout std_logic_vector(7 downto 0)  := (others => '0'); --   porta_a.export
		porta_b_export   : inout std_logic_vector(7 downto 0)  := (others => '0'); --   porta_b.export
		reset_reset_n    : in    std_logic                     := '0';             --     reset.reset_n
		saida_c_export   : out   std_logic_vector(7 downto 0);                     --   saida_c.export
		spi_MISO         : in    std_logic                     := '0';             --       spi.MISO
		spi_MOSI         : out   std_logic;                                        --          .MOSI
		spi_SCLK         : out   std_logic;                                        --          .SCLK
		spi_SS_n         : out   std_logic_vector(1 downto 0);                     --          .SS_n
		sw_export        : in    std_logic_vector(9 downto 0)  := (others => '0'); --        sw.export
		to_export        : out   std_logic;                                        --        to.export
		uart_rxd         : in    std_logic                     := '0';             --      uart.rxd
		uart_txd         : out   std_logic                                         --          .txd
	);
end entity sopc_2;

architecture rtl of sopc_2 is
	component sopc_2_PORTA_A is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component sopc_2_PORTA_A;

	component sopc_2_PORTA_B is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			irq        : out   std_logic                                         -- irq
		);
	end component sopc_2_PORTA_B;

	component sopc_2_botao is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component sopc_2_botao;

	component sopc_2_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component sopc_2_cpu;

	component sopc_2_entrada_C is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component sopc_2_entrada_C;

	component sopc_2_hex_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component sopc_2_hex_0;

	component sopc_2_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component sopc_2_jtag_uart;

	component sopc_2_memoria is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component sopc_2_memoria;

	component sopc_2_motor1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(13 downto 0)                     -- export
		);
	end component sopc_2_motor1;

	component sopc_2_saida_C is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component sopc_2_saida_C;

	component sopc_2_spi is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic_vector(1 downto 0)                      -- export
		);
	end component sopc_2_spi;

	component sopc_2_sw is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component sopc_2_sw;

	component sopc_2_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component sopc_2_sys_clk_timer;

	component sopc_2_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component sopc_2_sysid;

	component sopc_2_timer_geral is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			timeout_pulse : out std_logic                                         -- export
		);
	end component sopc_2_timer_geral;

	component sopc_2_timestamp_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component sopc_2_timestamp_timer;

	component sopc_2_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component sopc_2_uart;

	component sopc_2_watchdog_timer is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata     : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect   : in  std_logic                     := 'X';             -- chipselect
			write_n      : in  std_logic                     := 'X';             -- write_n
			irq          : out std_logic;                                        -- irq
			resetrequest : out std_logic                                         -- reset
		);
	end component sopc_2_watchdog_timer;

	component sopc_2_mm_interconnect_0 is
		port (
			clk_clk_clk                             : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                 : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			botao_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			botao_s1_write                          : out std_logic;                                        -- write
			botao_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			botao_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			botao_s1_chipselect                     : out std_logic;                                        -- chipselect
			cpu_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			entrada_C_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			entrada_C_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_0_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_0_s1_write                          : out std_logic;                                        -- write
			hex_0_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_0_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_1_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_1_s1_write                          : out std_logic;                                        -- write
			hex_1_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_1_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_1_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_2_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_2_s1_write                          : out std_logic;                                        -- write
			hex_2_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_2_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_2_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_3_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_3_s1_write                          : out std_logic;                                        -- write
			hex_3_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_3_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_3_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_4_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_4_s1_write                          : out std_logic;                                        -- write
			hex_4_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_4_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_4_s1_chipselect                     : out std_logic;                                        -- chipselect
			hex_5_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			hex_5_s1_write                          : out std_logic;                                        -- write
			hex_5_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_5_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			hex_5_s1_chipselect                     : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			memoria_s1_address                      : out std_logic_vector(13 downto 0);                    -- address
			memoria_s1_write                        : out std_logic;                                        -- write
			memoria_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			memoria_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			memoria_s1_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			memoria_s1_chipselect                   : out std_logic;                                        -- chipselect
			memoria_s1_clken                        : out std_logic;                                        -- clken
			motor1_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			motor1_s1_write                         : out std_logic;                                        -- write
			motor1_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			motor1_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			motor1_s1_chipselect                    : out std_logic;                                        -- chipselect
			motor2_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			motor2_s1_write                         : out std_logic;                                        -- write
			motor2_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			motor2_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			motor2_s1_chipselect                    : out std_logic;                                        -- chipselect
			motor3_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			motor3_s1_write                         : out std_logic;                                        -- write
			motor3_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			motor3_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			motor3_s1_chipselect                    : out std_logic;                                        -- chipselect
			motor4_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			motor4_s1_write                         : out std_logic;                                        -- write
			motor4_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			motor4_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			motor4_s1_chipselect                    : out std_logic;                                        -- chipselect
			PORTA_A_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			PORTA_A_s1_write                        : out std_logic;                                        -- write
			PORTA_A_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PORTA_A_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			PORTA_A_s1_chipselect                   : out std_logic;                                        -- chipselect
			PORTA_B_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			PORTA_B_s1_write                        : out std_logic;                                        -- write
			PORTA_B_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PORTA_B_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			PORTA_B_s1_chipselect                   : out std_logic;                                        -- chipselect
			saida_C_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			saida_C_s1_write                        : out std_logic;                                        -- write
			saida_C_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			saida_C_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			saida_C_s1_chipselect                   : out std_logic;                                        -- chipselect
			spi_spi_control_port_address            : out std_logic_vector(2 downto 0);                     -- address
			spi_spi_control_port_write              : out std_logic;                                        -- write
			spi_spi_control_port_read               : out std_logic;                                        -- read
			spi_spi_control_port_readdata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_spi_control_port_writedata          : out std_logic_vector(15 downto 0);                    -- writedata
			spi_spi_control_port_chipselect         : out std_logic;                                        -- chipselect
			sw_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			sw_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_address                : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                  : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata              : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect             : out std_logic;                                        -- chipselect
			sysid_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_geral_s1_address                  : out std_logic_vector(2 downto 0);                     -- address
			timer_geral_s1_write                    : out std_logic;                                        -- write
			timer_geral_s1_readdata                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_geral_s1_writedata                : out std_logic_vector(15 downto 0);                    -- writedata
			timer_geral_s1_chipselect               : out std_logic;                                        -- chipselect
			timestamp_timer_s1_address              : out std_logic_vector(2 downto 0);                     -- address
			timestamp_timer_s1_write                : out std_logic;                                        -- write
			timestamp_timer_s1_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timestamp_timer_s1_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			timestamp_timer_s1_chipselect           : out std_logic;                                        -- chipselect
			uart_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			uart_s1_write                           : out std_logic;                                        -- write
			uart_s1_read                            : out std_logic;                                        -- read
			uart_s1_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_s1_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			uart_s1_begintransfer                   : out std_logic;                                        -- begintransfer
			uart_s1_chipselect                      : out std_logic;                                        -- chipselect
			watchdog_timer_s1_address               : out std_logic_vector(2 downto 0);                     -- address
			watchdog_timer_s1_write                 : out std_logic;                                        -- write
			watchdog_timer_s1_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			watchdog_timer_s1_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			watchdog_timer_s1_chipselect            : out std_logic                                         -- chipselect
		);
	end component sopc_2_mm_interconnect_0;

	component sopc_2_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			receiver8_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component sopc_2_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                       : std_logic_vector(17 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(17 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest             : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_memoria_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:memoria_s1_chipselect -> memoria:chipselect
	signal mm_interconnect_0_memoria_s1_readdata                         : std_logic_vector(31 downto 0); -- memoria:readdata -> mm_interconnect_0:memoria_s1_readdata
	signal mm_interconnect_0_memoria_s1_address                          : std_logic_vector(13 downto 0); -- mm_interconnect_0:memoria_s1_address -> memoria:address
	signal mm_interconnect_0_memoria_s1_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:memoria_s1_byteenable -> memoria:byteenable
	signal mm_interconnect_0_memoria_s1_write                            : std_logic;                     -- mm_interconnect_0:memoria_s1_write -> memoria:write
	signal mm_interconnect_0_memoria_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:memoria_s1_writedata -> memoria:writedata
	signal mm_interconnect_0_memoria_s1_clken                            : std_logic;                     -- mm_interconnect_0:memoria_s1_clken -> memoria:clken
	signal mm_interconnect_0_porta_a_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:PORTA_A_s1_chipselect -> PORTA_A:chipselect
	signal mm_interconnect_0_porta_a_s1_readdata                         : std_logic_vector(31 downto 0); -- PORTA_A:readdata -> mm_interconnect_0:PORTA_A_s1_readdata
	signal mm_interconnect_0_porta_a_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:PORTA_A_s1_address -> PORTA_A:address
	signal mm_interconnect_0_porta_a_s1_write                            : std_logic;                     -- mm_interconnect_0:PORTA_A_s1_write -> mm_interconnect_0_porta_a_s1_write:in
	signal mm_interconnect_0_porta_a_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:PORTA_A_s1_writedata -> PORTA_A:writedata
	signal mm_interconnect_0_porta_b_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:PORTA_B_s1_chipselect -> PORTA_B:chipselect
	signal mm_interconnect_0_porta_b_s1_readdata                         : std_logic_vector(31 downto 0); -- PORTA_B:readdata -> mm_interconnect_0:PORTA_B_s1_readdata
	signal mm_interconnect_0_porta_b_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:PORTA_B_s1_address -> PORTA_B:address
	signal mm_interconnect_0_porta_b_s1_write                            : std_logic;                     -- mm_interconnect_0:PORTA_B_s1_write -> mm_interconnect_0_porta_b_s1_write:in
	signal mm_interconnect_0_porta_b_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:PORTA_B_s1_writedata -> PORTA_B:writedata
	signal mm_interconnect_0_saida_c_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:saida_C_s1_chipselect -> saida_C:chipselect
	signal mm_interconnect_0_saida_c_s1_readdata                         : std_logic_vector(31 downto 0); -- saida_C:readdata -> mm_interconnect_0:saida_C_s1_readdata
	signal mm_interconnect_0_saida_c_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:saida_C_s1_address -> saida_C:address
	signal mm_interconnect_0_saida_c_s1_write                            : std_logic;                     -- mm_interconnect_0:saida_C_s1_write -> mm_interconnect_0_saida_c_s1_write:in
	signal mm_interconnect_0_saida_c_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:saida_C_s1_writedata -> saida_C:writedata
	signal mm_interconnect_0_entrada_c_s1_readdata                       : std_logic_vector(31 downto 0); -- entrada_C:readdata -> mm_interconnect_0:entrada_C_s1_readdata
	signal mm_interconnect_0_entrada_c_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:entrada_C_s1_address -> entrada_C:address
	signal mm_interconnect_0_uart_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                            : std_logic_vector(15 downto 0); -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                                : std_logic;                     -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer                       : std_logic;                     -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                               : std_logic;                     -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal mm_interconnect_0_botao_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:botao_s1_chipselect -> botao:chipselect
	signal mm_interconnect_0_botao_s1_readdata                           : std_logic_vector(31 downto 0); -- botao:readdata -> mm_interconnect_0:botao_s1_readdata
	signal mm_interconnect_0_botao_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:botao_s1_address -> botao:address
	signal mm_interconnect_0_botao_s1_write                              : std_logic;                     -- mm_interconnect_0:botao_s1_write -> mm_interconnect_0_botao_s1_write:in
	signal mm_interconnect_0_botao_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:botao_s1_writedata -> botao:writedata
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                   : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                      : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_timestamp_timer_s1_chipselect               : std_logic;                     -- mm_interconnect_0:timestamp_timer_s1_chipselect -> timestamp_timer:chipselect
	signal mm_interconnect_0_timestamp_timer_s1_readdata                 : std_logic_vector(15 downto 0); -- timestamp_timer:readdata -> mm_interconnect_0:timestamp_timer_s1_readdata
	signal mm_interconnect_0_timestamp_timer_s1_address                  : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timestamp_timer_s1_address -> timestamp_timer:address
	signal mm_interconnect_0_timestamp_timer_s1_write                    : std_logic;                     -- mm_interconnect_0:timestamp_timer_s1_write -> mm_interconnect_0_timestamp_timer_s1_write:in
	signal mm_interconnect_0_timestamp_timer_s1_writedata                : std_logic_vector(15 downto 0); -- mm_interconnect_0:timestamp_timer_s1_writedata -> timestamp_timer:writedata
	signal mm_interconnect_0_timer_geral_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:timer_geral_s1_chipselect -> timer_geral:chipselect
	signal mm_interconnect_0_timer_geral_s1_readdata                     : std_logic_vector(15 downto 0); -- timer_geral:readdata -> mm_interconnect_0:timer_geral_s1_readdata
	signal mm_interconnect_0_timer_geral_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_geral_s1_address -> timer_geral:address
	signal mm_interconnect_0_timer_geral_s1_write                        : std_logic;                     -- mm_interconnect_0:timer_geral_s1_write -> mm_interconnect_0_timer_geral_s1_write:in
	signal mm_interconnect_0_timer_geral_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_geral_s1_writedata -> timer_geral:writedata
	signal mm_interconnect_0_watchdog_timer_s1_chipselect                : std_logic;                     -- mm_interconnect_0:watchdog_timer_s1_chipselect -> watchdog_timer:chipselect
	signal mm_interconnect_0_watchdog_timer_s1_readdata                  : std_logic_vector(15 downto 0); -- watchdog_timer:readdata -> mm_interconnect_0:watchdog_timer_s1_readdata
	signal mm_interconnect_0_watchdog_timer_s1_address                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:watchdog_timer_s1_address -> watchdog_timer:address
	signal mm_interconnect_0_watchdog_timer_s1_write                     : std_logic;                     -- mm_interconnect_0:watchdog_timer_s1_write -> mm_interconnect_0_watchdog_timer_s1_write:in
	signal mm_interconnect_0_watchdog_timer_s1_writedata                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:watchdog_timer_s1_writedata -> watchdog_timer:writedata
	signal mm_interconnect_0_hex_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:hex_0_s1_chipselect -> hex_0:chipselect
	signal mm_interconnect_0_hex_0_s1_readdata                           : std_logic_vector(31 downto 0); -- hex_0:readdata -> mm_interconnect_0:hex_0_s1_readdata
	signal mm_interconnect_0_hex_0_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_0_s1_address -> hex_0:address
	signal mm_interconnect_0_hex_0_s1_write                              : std_logic;                     -- mm_interconnect_0:hex_0_s1_write -> mm_interconnect_0_hex_0_s1_write:in
	signal mm_interconnect_0_hex_0_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_0_s1_writedata -> hex_0:writedata
	signal mm_interconnect_0_hex_5_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:hex_5_s1_chipselect -> hex_5:chipselect
	signal mm_interconnect_0_hex_5_s1_readdata                           : std_logic_vector(31 downto 0); -- hex_5:readdata -> mm_interconnect_0:hex_5_s1_readdata
	signal mm_interconnect_0_hex_5_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_5_s1_address -> hex_5:address
	signal mm_interconnect_0_hex_5_s1_write                              : std_logic;                     -- mm_interconnect_0:hex_5_s1_write -> mm_interconnect_0_hex_5_s1_write:in
	signal mm_interconnect_0_hex_5_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_5_s1_writedata -> hex_5:writedata
	signal mm_interconnect_0_hex_4_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:hex_4_s1_chipselect -> hex_4:chipselect
	signal mm_interconnect_0_hex_4_s1_readdata                           : std_logic_vector(31 downto 0); -- hex_4:readdata -> mm_interconnect_0:hex_4_s1_readdata
	signal mm_interconnect_0_hex_4_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_4_s1_address -> hex_4:address
	signal mm_interconnect_0_hex_4_s1_write                              : std_logic;                     -- mm_interconnect_0:hex_4_s1_write -> mm_interconnect_0_hex_4_s1_write:in
	signal mm_interconnect_0_hex_4_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_4_s1_writedata -> hex_4:writedata
	signal mm_interconnect_0_hex_3_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:hex_3_s1_chipselect -> hex_3:chipselect
	signal mm_interconnect_0_hex_3_s1_readdata                           : std_logic_vector(31 downto 0); -- hex_3:readdata -> mm_interconnect_0:hex_3_s1_readdata
	signal mm_interconnect_0_hex_3_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_3_s1_address -> hex_3:address
	signal mm_interconnect_0_hex_3_s1_write                              : std_logic;                     -- mm_interconnect_0:hex_3_s1_write -> mm_interconnect_0_hex_3_s1_write:in
	signal mm_interconnect_0_hex_3_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_3_s1_writedata -> hex_3:writedata
	signal mm_interconnect_0_hex_2_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:hex_2_s1_chipselect -> hex_2:chipselect
	signal mm_interconnect_0_hex_2_s1_readdata                           : std_logic_vector(31 downto 0); -- hex_2:readdata -> mm_interconnect_0:hex_2_s1_readdata
	signal mm_interconnect_0_hex_2_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_2_s1_address -> hex_2:address
	signal mm_interconnect_0_hex_2_s1_write                              : std_logic;                     -- mm_interconnect_0:hex_2_s1_write -> mm_interconnect_0_hex_2_s1_write:in
	signal mm_interconnect_0_hex_2_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_2_s1_writedata -> hex_2:writedata
	signal mm_interconnect_0_hex_1_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:hex_1_s1_chipselect -> hex_1:chipselect
	signal mm_interconnect_0_hex_1_s1_readdata                           : std_logic_vector(31 downto 0); -- hex_1:readdata -> mm_interconnect_0:hex_1_s1_readdata
	signal mm_interconnect_0_hex_1_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_1_s1_address -> hex_1:address
	signal mm_interconnect_0_hex_1_s1_write                              : std_logic;                     -- mm_interconnect_0:hex_1_s1_write -> mm_interconnect_0_hex_1_s1_write:in
	signal mm_interconnect_0_hex_1_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_1_s1_writedata -> hex_1:writedata
	signal mm_interconnect_0_sw_s1_readdata                              : std_logic_vector(31 downto 0); -- sw:readdata -> mm_interconnect_0:sw_s1_readdata
	signal mm_interconnect_0_sw_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sw_s1_address -> sw:address
	signal mm_interconnect_0_motor1_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:motor1_s1_chipselect -> motor1:chipselect
	signal mm_interconnect_0_motor1_s1_readdata                          : std_logic_vector(31 downto 0); -- motor1:readdata -> mm_interconnect_0:motor1_s1_readdata
	signal mm_interconnect_0_motor1_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:motor1_s1_address -> motor1:address
	signal mm_interconnect_0_motor1_s1_write                             : std_logic;                     -- mm_interconnect_0:motor1_s1_write -> mm_interconnect_0_motor1_s1_write:in
	signal mm_interconnect_0_motor1_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:motor1_s1_writedata -> motor1:writedata
	signal mm_interconnect_0_motor2_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:motor2_s1_chipselect -> motor2:chipselect
	signal mm_interconnect_0_motor2_s1_readdata                          : std_logic_vector(31 downto 0); -- motor2:readdata -> mm_interconnect_0:motor2_s1_readdata
	signal mm_interconnect_0_motor2_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:motor2_s1_address -> motor2:address
	signal mm_interconnect_0_motor2_s1_write                             : std_logic;                     -- mm_interconnect_0:motor2_s1_write -> mm_interconnect_0_motor2_s1_write:in
	signal mm_interconnect_0_motor2_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:motor2_s1_writedata -> motor2:writedata
	signal mm_interconnect_0_motor4_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:motor4_s1_chipselect -> motor4:chipselect
	signal mm_interconnect_0_motor4_s1_readdata                          : std_logic_vector(31 downto 0); -- motor4:readdata -> mm_interconnect_0:motor4_s1_readdata
	signal mm_interconnect_0_motor4_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:motor4_s1_address -> motor4:address
	signal mm_interconnect_0_motor4_s1_write                             : std_logic;                     -- mm_interconnect_0:motor4_s1_write -> mm_interconnect_0_motor4_s1_write:in
	signal mm_interconnect_0_motor4_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:motor4_s1_writedata -> motor4:writedata
	signal mm_interconnect_0_motor3_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:motor3_s1_chipselect -> motor3:chipselect
	signal mm_interconnect_0_motor3_s1_readdata                          : std_logic_vector(31 downto 0); -- motor3:readdata -> mm_interconnect_0:motor3_s1_readdata
	signal mm_interconnect_0_motor3_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:motor3_s1_address -> motor3:address
	signal mm_interconnect_0_motor3_s1_write                             : std_logic;                     -- mm_interconnect_0:motor3_s1_write -> mm_interconnect_0_motor3_s1_write:in
	signal mm_interconnect_0_motor3_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:motor3_s1_writedata -> motor3:writedata
	signal mm_interconnect_0_spi_spi_control_port_chipselect             : std_logic;                     -- mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	signal mm_interconnect_0_spi_spi_control_port_readdata               : std_logic_vector(15 downto 0); -- spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	signal mm_interconnect_0_spi_spi_control_port_address                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	signal mm_interconnect_0_spi_spi_control_port_read                   : std_logic;                     -- mm_interconnect_0:spi_spi_control_port_read -> mm_interconnect_0_spi_spi_control_port_read:in
	signal mm_interconnect_0_spi_spi_control_port_write                  : std_logic;                     -- mm_interconnect_0:spi_spi_control_port_write -> mm_interconnect_0_spi_spi_control_port_write:in
	signal mm_interconnect_0_spi_spi_control_port_writedata              : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- PORTA_B:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- uart:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- spi:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                      : std_logic;                     -- botao:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                      : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                      : std_logic;                     -- timestamp_timer:irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                      : std_logic;                     -- timer_geral:irq -> irq_mapper:receiver7_irq
	signal irq_mapper_receiver8_irq                                      : std_logic;                     -- watchdog_timer:irq -> irq_mapper:receiver8_irq
	signal cpu_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, memoria:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, memoria:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                 : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in1
	signal watchdog_timer_resetrequest_reset                             : std_logic;                     -- watchdog_timer:resetrequest -> rst_controller:reset_in2
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_porta_a_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_porta_a_s1_write:inv -> PORTA_A:write_n
	signal mm_interconnect_0_porta_b_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_porta_b_s1_write:inv -> PORTA_B:write_n
	signal mm_interconnect_0_saida_c_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_saida_c_s1_write:inv -> saida_C:write_n
	signal mm_interconnect_0_uart_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal mm_interconnect_0_botao_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_botao_s1_write:inv -> botao:write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_0_timestamp_timer_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_0_timestamp_timer_s1_write:inv -> timestamp_timer:write_n
	signal mm_interconnect_0_timer_geral_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_timer_geral_s1_write:inv -> timer_geral:write_n
	signal mm_interconnect_0_watchdog_timer_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_watchdog_timer_s1_write:inv -> watchdog_timer:write_n
	signal mm_interconnect_0_hex_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_hex_0_s1_write:inv -> hex_0:write_n
	signal mm_interconnect_0_hex_5_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_hex_5_s1_write:inv -> hex_5:write_n
	signal mm_interconnect_0_hex_4_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_hex_4_s1_write:inv -> hex_4:write_n
	signal mm_interconnect_0_hex_3_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_hex_3_s1_write:inv -> hex_3:write_n
	signal mm_interconnect_0_hex_2_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_hex_2_s1_write:inv -> hex_2:write_n
	signal mm_interconnect_0_hex_1_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_hex_1_s1_write:inv -> hex_1:write_n
	signal mm_interconnect_0_motor1_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_motor1_s1_write:inv -> motor1:write_n
	signal mm_interconnect_0_motor2_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_motor2_s1_write:inv -> motor2:write_n
	signal mm_interconnect_0_motor4_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_motor4_s1_write:inv -> motor4:write_n
	signal mm_interconnect_0_motor3_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_motor3_s1_write:inv -> motor3:write_n
	signal mm_interconnect_0_spi_spi_control_port_read_ports_inv         : std_logic;                     -- mm_interconnect_0_spi_spi_control_port_read:inv -> spi:read_n
	signal mm_interconnect_0_spi_spi_control_port_write_ports_inv        : std_logic;                     -- mm_interconnect_0_spi_spi_control_port_write:inv -> spi:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [PORTA_A:reset_n, PORTA_B:reset_n, botao:reset_n, cpu:reset_n, entrada_C:reset_n, hex_0:reset_n, hex_1:reset_n, hex_2:reset_n, hex_3:reset_n, hex_4:reset_n, hex_5:reset_n, jtag_uart:rst_n, motor1:reset_n, motor2:reset_n, motor3:reset_n, motor4:reset_n, saida_C:reset_n, spi:reset_n, sw:reset_n, sys_clk_timer:reset_n, sysid:reset_n, timer_geral:reset_n, timestamp_timer:reset_n, uart:reset_n, watchdog_timer:reset_n]

begin

	porta_a : component sopc_2_PORTA_A
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_porta_a_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_porta_a_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_porta_a_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_porta_a_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_porta_a_s1_readdata,        --                    .readdata
			bidir_port => porta_a_export                                -- external_connection.export
		);

	porta_b : component sopc_2_PORTA_B
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_porta_b_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_porta_b_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_porta_b_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_porta_b_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_porta_b_s1_readdata,        --                    .readdata
			bidir_port => porta_b_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                      --                 irq.irq
		);

	botao : component sopc_2_botao
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_botao_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_botao_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_botao_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_botao_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_botao_s1_readdata,        --                    .readdata
			in_port    => botao_export,                               -- external_connection.export
			irq        => irq_mapper_receiver4_irq                    --                 irq.irq
		);

	cpu : component sopc_2_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	entrada_c : component sopc_2_entrada_C
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_entrada_c_s1_address,   --                  s1.address
			readdata => mm_interconnect_0_entrada_c_s1_readdata,  --                    .readdata
			in_port  => entrada_c_export                          -- external_connection.export
		);

	hex_0 : component sopc_2_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_0_s1_readdata,        --                    .readdata
			out_port   => hex0_export                                 -- external_connection.export
		);

	hex_1 : component sopc_2_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_1_s1_readdata,        --                    .readdata
			out_port   => hex1_export                                 -- external_connection.export
		);

	hex_2 : component sopc_2_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_2_s1_readdata,        --                    .readdata
			out_port   => hex2_export                                 -- external_connection.export
		);

	hex_3 : component sopc_2_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_3_s1_readdata,        --                    .readdata
			out_port   => hex3_export                                 -- external_connection.export
		);

	hex_4 : component sopc_2_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_4_s1_readdata,        --                    .readdata
			out_port   => hex_4_export                                -- external_connection.export
		);

	hex_5 : component sopc_2_hex_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_hex_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_5_s1_readdata,        --                    .readdata
			out_port   => hex5_export                                 -- external_connection.export
		);

	jtag_uart : component sopc_2_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	memoria : component sopc_2_memoria
		port map (
			clk        => clk_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_memoria_s1_address,    --     s1.address
			clken      => mm_interconnect_0_memoria_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_memoria_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_memoria_s1_write,      --       .write
			readdata   => mm_interconnect_0_memoria_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_memoria_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_memoria_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,          -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,      --       .reset_req
			freeze     => '0'                                      -- (terminated)
		);

	motor1 : component sopc_2_motor1
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_motor1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motor1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motor1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motor1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motor1_s1_readdata,        --                    .readdata
			out_port   => motor_1_export                               -- external_connection.export
		);

	motor2 : component sopc_2_motor1
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_motor2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motor2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motor2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motor2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motor2_s1_readdata,        --                    .readdata
			out_port   => motor2_export                                -- external_connection.export
		);

	motor3 : component sopc_2_motor1
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_motor3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motor3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motor3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motor3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motor3_s1_readdata,        --                    .readdata
			out_port   => motor3_export                                -- external_connection.export
		);

	motor4 : component sopc_2_motor1
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_motor4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motor4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motor4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motor4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motor4_s1_readdata,        --                    .readdata
			out_port   => motor4_export                                -- external_connection.export
		);

	saida_c : component sopc_2_saida_C
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_saida_c_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_saida_c_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_saida_c_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_saida_c_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_saida_c_s1_readdata,        --                    .readdata
			out_port   => saida_c_export                                -- external_connection.export
		);

	spi : component sopc_2_spi
		port map (
			clk           => clk_clk,                                                --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,               --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver3_irq,                               --              irq.irq
			MISO          => spi_MISO,                                               --         external.export
			MOSI          => spi_MOSI,                                               --                 .export
			SCLK          => spi_SCLK,                                               --                 .export
			SS_n          => spi_SS_n                                                --                 .export
		);

	sw : component sopc_2_sw
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_sw_s1_address,          --                  s1.address
			readdata => mm_interconnect_0_sw_s1_readdata,         --                    .readdata
			in_port  => sw_export                                 -- external_connection.export
		);

	sys_clk_timer : component sopc_2_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver5_irq                            --   irq.irq
		);

	sysid : component sopc_2_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer_geral : component sopc_2_timer_geral
		port map (
			clk           => clk_clk,                                          --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			address       => mm_interconnect_0_timer_geral_s1_address,         --            s1.address
			writedata     => mm_interconnect_0_timer_geral_s1_writedata,       --              .writedata
			readdata      => mm_interconnect_0_timer_geral_s1_readdata,        --              .readdata
			chipselect    => mm_interconnect_0_timer_geral_s1_chipselect,      --              .chipselect
			write_n       => mm_interconnect_0_timer_geral_s1_write_ports_inv, --              .write_n
			irq           => irq_mapper_receiver7_irq,                         --           irq.irq
			timeout_pulse => to_export                                         -- external_port.export
		);

	timestamp_timer : component sopc_2_timestamp_timer
		port map (
			clk        => clk_clk,                                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             -- reset.reset_n
			address    => mm_interconnect_0_timestamp_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timestamp_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timestamp_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timestamp_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timestamp_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver6_irq                              --   irq.irq
		);

	uart : component sopc_2_uart
		port map (
			clk           => clk_clk,                                   --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			rxd           => uart_rxd,                                  -- external_connection.export
			txd           => uart_txd,                                  --                    .export
			irq           => irq_mapper_receiver2_irq                   --                 irq.irq
		);

	watchdog_timer : component sopc_2_watchdog_timer
		port map (
			clk          => clk_clk,                                             --          clk.clk
			reset_n      => rst_controller_reset_out_reset_ports_inv,            --        reset.reset_n
			address      => mm_interconnect_0_watchdog_timer_s1_address,         --           s1.address
			writedata    => mm_interconnect_0_watchdog_timer_s1_writedata,       --             .writedata
			readdata     => mm_interconnect_0_watchdog_timer_s1_readdata,        --             .readdata
			chipselect   => mm_interconnect_0_watchdog_timer_s1_chipselect,      --             .chipselect
			write_n      => mm_interconnect_0_watchdog_timer_s1_write_ports_inv, --             .write_n
			irq          => irq_mapper_receiver8_irq,                            --          irq.irq
			resetrequest => watchdog_timer_resetrequest_reset                    -- resetrequest.reset
		);

	mm_interconnect_0 : component sopc_2_mm_interconnect_0
		port map (
			clk_clk_clk                             => clk_clk,                                                   --                         clk_clk.clk
			cpu_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                            -- cpu_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                 => cpu_data_master_address,                                   --                 cpu_data_master.address
			cpu_data_master_waitrequest             => cpu_data_master_waitrequest,                               --                                .waitrequest
			cpu_data_master_byteenable              => cpu_data_master_byteenable,                                --                                .byteenable
			cpu_data_master_read                    => cpu_data_master_read,                                      --                                .read
			cpu_data_master_readdata                => cpu_data_master_readdata,                                  --                                .readdata
			cpu_data_master_write                   => cpu_data_master_write,                                     --                                .write
			cpu_data_master_writedata               => cpu_data_master_writedata,                                 --                                .writedata
			cpu_data_master_debugaccess             => cpu_data_master_debugaccess,                               --                                .debugaccess
			cpu_instruction_master_address          => cpu_instruction_master_address,                            --          cpu_instruction_master.address
			cpu_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                        --                                .waitrequest
			cpu_instruction_master_read             => cpu_instruction_master_read,                               --                                .read
			cpu_instruction_master_readdata         => cpu_instruction_master_readdata,                           --                                .readdata
			botao_s1_address                        => mm_interconnect_0_botao_s1_address,                        --                        botao_s1.address
			botao_s1_write                          => mm_interconnect_0_botao_s1_write,                          --                                .write
			botao_s1_readdata                       => mm_interconnect_0_botao_s1_readdata,                       --                                .readdata
			botao_s1_writedata                      => mm_interconnect_0_botao_s1_writedata,                      --                                .writedata
			botao_s1_chipselect                     => mm_interconnect_0_botao_s1_chipselect,                     --                                .chipselect
			cpu_debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,             --             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                .write
			cpu_debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                .read
			cpu_debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                .readdata
			cpu_debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                .writedata
			cpu_debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                .byteenable
			cpu_debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                .waitrequest
			cpu_debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                .debugaccess
			entrada_C_s1_address                    => mm_interconnect_0_entrada_c_s1_address,                    --                    entrada_C_s1.address
			entrada_C_s1_readdata                   => mm_interconnect_0_entrada_c_s1_readdata,                   --                                .readdata
			hex_0_s1_address                        => mm_interconnect_0_hex_0_s1_address,                        --                        hex_0_s1.address
			hex_0_s1_write                          => mm_interconnect_0_hex_0_s1_write,                          --                                .write
			hex_0_s1_readdata                       => mm_interconnect_0_hex_0_s1_readdata,                       --                                .readdata
			hex_0_s1_writedata                      => mm_interconnect_0_hex_0_s1_writedata,                      --                                .writedata
			hex_0_s1_chipselect                     => mm_interconnect_0_hex_0_s1_chipselect,                     --                                .chipselect
			hex_1_s1_address                        => mm_interconnect_0_hex_1_s1_address,                        --                        hex_1_s1.address
			hex_1_s1_write                          => mm_interconnect_0_hex_1_s1_write,                          --                                .write
			hex_1_s1_readdata                       => mm_interconnect_0_hex_1_s1_readdata,                       --                                .readdata
			hex_1_s1_writedata                      => mm_interconnect_0_hex_1_s1_writedata,                      --                                .writedata
			hex_1_s1_chipselect                     => mm_interconnect_0_hex_1_s1_chipselect,                     --                                .chipselect
			hex_2_s1_address                        => mm_interconnect_0_hex_2_s1_address,                        --                        hex_2_s1.address
			hex_2_s1_write                          => mm_interconnect_0_hex_2_s1_write,                          --                                .write
			hex_2_s1_readdata                       => mm_interconnect_0_hex_2_s1_readdata,                       --                                .readdata
			hex_2_s1_writedata                      => mm_interconnect_0_hex_2_s1_writedata,                      --                                .writedata
			hex_2_s1_chipselect                     => mm_interconnect_0_hex_2_s1_chipselect,                     --                                .chipselect
			hex_3_s1_address                        => mm_interconnect_0_hex_3_s1_address,                        --                        hex_3_s1.address
			hex_3_s1_write                          => mm_interconnect_0_hex_3_s1_write,                          --                                .write
			hex_3_s1_readdata                       => mm_interconnect_0_hex_3_s1_readdata,                       --                                .readdata
			hex_3_s1_writedata                      => mm_interconnect_0_hex_3_s1_writedata,                      --                                .writedata
			hex_3_s1_chipselect                     => mm_interconnect_0_hex_3_s1_chipselect,                     --                                .chipselect
			hex_4_s1_address                        => mm_interconnect_0_hex_4_s1_address,                        --                        hex_4_s1.address
			hex_4_s1_write                          => mm_interconnect_0_hex_4_s1_write,                          --                                .write
			hex_4_s1_readdata                       => mm_interconnect_0_hex_4_s1_readdata,                       --                                .readdata
			hex_4_s1_writedata                      => mm_interconnect_0_hex_4_s1_writedata,                      --                                .writedata
			hex_4_s1_chipselect                     => mm_interconnect_0_hex_4_s1_chipselect,                     --                                .chipselect
			hex_5_s1_address                        => mm_interconnect_0_hex_5_s1_address,                        --                        hex_5_s1.address
			hex_5_s1_write                          => mm_interconnect_0_hex_5_s1_write,                          --                                .write
			hex_5_s1_readdata                       => mm_interconnect_0_hex_5_s1_readdata,                       --                                .readdata
			hex_5_s1_writedata                      => mm_interconnect_0_hex_5_s1_writedata,                      --                                .writedata
			hex_5_s1_chipselect                     => mm_interconnect_0_hex_5_s1_chipselect,                     --                                .chipselect
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                .chipselect
			memoria_s1_address                      => mm_interconnect_0_memoria_s1_address,                      --                      memoria_s1.address
			memoria_s1_write                        => mm_interconnect_0_memoria_s1_write,                        --                                .write
			memoria_s1_readdata                     => mm_interconnect_0_memoria_s1_readdata,                     --                                .readdata
			memoria_s1_writedata                    => mm_interconnect_0_memoria_s1_writedata,                    --                                .writedata
			memoria_s1_byteenable                   => mm_interconnect_0_memoria_s1_byteenable,                   --                                .byteenable
			memoria_s1_chipselect                   => mm_interconnect_0_memoria_s1_chipselect,                   --                                .chipselect
			memoria_s1_clken                        => mm_interconnect_0_memoria_s1_clken,                        --                                .clken
			motor1_s1_address                       => mm_interconnect_0_motor1_s1_address,                       --                       motor1_s1.address
			motor1_s1_write                         => mm_interconnect_0_motor1_s1_write,                         --                                .write
			motor1_s1_readdata                      => mm_interconnect_0_motor1_s1_readdata,                      --                                .readdata
			motor1_s1_writedata                     => mm_interconnect_0_motor1_s1_writedata,                     --                                .writedata
			motor1_s1_chipselect                    => mm_interconnect_0_motor1_s1_chipselect,                    --                                .chipselect
			motor2_s1_address                       => mm_interconnect_0_motor2_s1_address,                       --                       motor2_s1.address
			motor2_s1_write                         => mm_interconnect_0_motor2_s1_write,                         --                                .write
			motor2_s1_readdata                      => mm_interconnect_0_motor2_s1_readdata,                      --                                .readdata
			motor2_s1_writedata                     => mm_interconnect_0_motor2_s1_writedata,                     --                                .writedata
			motor2_s1_chipselect                    => mm_interconnect_0_motor2_s1_chipselect,                    --                                .chipselect
			motor3_s1_address                       => mm_interconnect_0_motor3_s1_address,                       --                       motor3_s1.address
			motor3_s1_write                         => mm_interconnect_0_motor3_s1_write,                         --                                .write
			motor3_s1_readdata                      => mm_interconnect_0_motor3_s1_readdata,                      --                                .readdata
			motor3_s1_writedata                     => mm_interconnect_0_motor3_s1_writedata,                     --                                .writedata
			motor3_s1_chipselect                    => mm_interconnect_0_motor3_s1_chipselect,                    --                                .chipselect
			motor4_s1_address                       => mm_interconnect_0_motor4_s1_address,                       --                       motor4_s1.address
			motor4_s1_write                         => mm_interconnect_0_motor4_s1_write,                         --                                .write
			motor4_s1_readdata                      => mm_interconnect_0_motor4_s1_readdata,                      --                                .readdata
			motor4_s1_writedata                     => mm_interconnect_0_motor4_s1_writedata,                     --                                .writedata
			motor4_s1_chipselect                    => mm_interconnect_0_motor4_s1_chipselect,                    --                                .chipselect
			PORTA_A_s1_address                      => mm_interconnect_0_porta_a_s1_address,                      --                      PORTA_A_s1.address
			PORTA_A_s1_write                        => mm_interconnect_0_porta_a_s1_write,                        --                                .write
			PORTA_A_s1_readdata                     => mm_interconnect_0_porta_a_s1_readdata,                     --                                .readdata
			PORTA_A_s1_writedata                    => mm_interconnect_0_porta_a_s1_writedata,                    --                                .writedata
			PORTA_A_s1_chipselect                   => mm_interconnect_0_porta_a_s1_chipselect,                   --                                .chipselect
			PORTA_B_s1_address                      => mm_interconnect_0_porta_b_s1_address,                      --                      PORTA_B_s1.address
			PORTA_B_s1_write                        => mm_interconnect_0_porta_b_s1_write,                        --                                .write
			PORTA_B_s1_readdata                     => mm_interconnect_0_porta_b_s1_readdata,                     --                                .readdata
			PORTA_B_s1_writedata                    => mm_interconnect_0_porta_b_s1_writedata,                    --                                .writedata
			PORTA_B_s1_chipselect                   => mm_interconnect_0_porta_b_s1_chipselect,                   --                                .chipselect
			saida_C_s1_address                      => mm_interconnect_0_saida_c_s1_address,                      --                      saida_C_s1.address
			saida_C_s1_write                        => mm_interconnect_0_saida_c_s1_write,                        --                                .write
			saida_C_s1_readdata                     => mm_interconnect_0_saida_c_s1_readdata,                     --                                .readdata
			saida_C_s1_writedata                    => mm_interconnect_0_saida_c_s1_writedata,                    --                                .writedata
			saida_C_s1_chipselect                   => mm_interconnect_0_saida_c_s1_chipselect,                   --                                .chipselect
			spi_spi_control_port_address            => mm_interconnect_0_spi_spi_control_port_address,            --            spi_spi_control_port.address
			spi_spi_control_port_write              => mm_interconnect_0_spi_spi_control_port_write,              --                                .write
			spi_spi_control_port_read               => mm_interconnect_0_spi_spi_control_port_read,               --                                .read
			spi_spi_control_port_readdata           => mm_interconnect_0_spi_spi_control_port_readdata,           --                                .readdata
			spi_spi_control_port_writedata          => mm_interconnect_0_spi_spi_control_port_writedata,          --                                .writedata
			spi_spi_control_port_chipselect         => mm_interconnect_0_spi_spi_control_port_chipselect,         --                                .chipselect
			sw_s1_address                           => mm_interconnect_0_sw_s1_address,                           --                           sw_s1.address
			sw_s1_readdata                          => mm_interconnect_0_sw_s1_readdata,                          --                                .readdata
			sys_clk_timer_s1_address                => mm_interconnect_0_sys_clk_timer_s1_address,                --                sys_clk_timer_s1.address
			sys_clk_timer_s1_write                  => mm_interconnect_0_sys_clk_timer_s1_write,                  --                                .write
			sys_clk_timer_s1_readdata               => mm_interconnect_0_sys_clk_timer_s1_readdata,               --                                .readdata
			sys_clk_timer_s1_writedata              => mm_interconnect_0_sys_clk_timer_s1_writedata,              --                                .writedata
			sys_clk_timer_s1_chipselect             => mm_interconnect_0_sys_clk_timer_s1_chipselect,             --                                .chipselect
			sysid_control_slave_address             => mm_interconnect_0_sysid_control_slave_address,             --             sysid_control_slave.address
			sysid_control_slave_readdata            => mm_interconnect_0_sysid_control_slave_readdata,            --                                .readdata
			timer_geral_s1_address                  => mm_interconnect_0_timer_geral_s1_address,                  --                  timer_geral_s1.address
			timer_geral_s1_write                    => mm_interconnect_0_timer_geral_s1_write,                    --                                .write
			timer_geral_s1_readdata                 => mm_interconnect_0_timer_geral_s1_readdata,                 --                                .readdata
			timer_geral_s1_writedata                => mm_interconnect_0_timer_geral_s1_writedata,                --                                .writedata
			timer_geral_s1_chipselect               => mm_interconnect_0_timer_geral_s1_chipselect,               --                                .chipselect
			timestamp_timer_s1_address              => mm_interconnect_0_timestamp_timer_s1_address,              --              timestamp_timer_s1.address
			timestamp_timer_s1_write                => mm_interconnect_0_timestamp_timer_s1_write,                --                                .write
			timestamp_timer_s1_readdata             => mm_interconnect_0_timestamp_timer_s1_readdata,             --                                .readdata
			timestamp_timer_s1_writedata            => mm_interconnect_0_timestamp_timer_s1_writedata,            --                                .writedata
			timestamp_timer_s1_chipselect           => mm_interconnect_0_timestamp_timer_s1_chipselect,           --                                .chipselect
			uart_s1_address                         => mm_interconnect_0_uart_s1_address,                         --                         uart_s1.address
			uart_s1_write                           => mm_interconnect_0_uart_s1_write,                           --                                .write
			uart_s1_read                            => mm_interconnect_0_uart_s1_read,                            --                                .read
			uart_s1_readdata                        => mm_interconnect_0_uart_s1_readdata,                        --                                .readdata
			uart_s1_writedata                       => mm_interconnect_0_uart_s1_writedata,                       --                                .writedata
			uart_s1_begintransfer                   => mm_interconnect_0_uart_s1_begintransfer,                   --                                .begintransfer
			uart_s1_chipselect                      => mm_interconnect_0_uart_s1_chipselect,                      --                                .chipselect
			watchdog_timer_s1_address               => mm_interconnect_0_watchdog_timer_s1_address,               --               watchdog_timer_s1.address
			watchdog_timer_s1_write                 => mm_interconnect_0_watchdog_timer_s1_write,                 --                                .write
			watchdog_timer_s1_readdata              => mm_interconnect_0_watchdog_timer_s1_readdata,              --                                .readdata
			watchdog_timer_s1_writedata             => mm_interconnect_0_watchdog_timer_s1_writedata,             --                                .writedata
			watchdog_timer_s1_chipselect            => mm_interconnect_0_watchdog_timer_s1_chipselect             --                                .chipselect
		);

	irq_mapper : component sopc_2_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,       -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,       -- receiver7.irq
			receiver8_irq => irq_mapper_receiver8_irq,       -- receiver8.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			reset_in2      => watchdog_timer_resetrequest_reset,  -- reset_in2.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_porta_a_s1_write_ports_inv <= not mm_interconnect_0_porta_a_s1_write;

	mm_interconnect_0_porta_b_s1_write_ports_inv <= not mm_interconnect_0_porta_b_s1_write;

	mm_interconnect_0_saida_c_s1_write_ports_inv <= not mm_interconnect_0_saida_c_s1_write;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	mm_interconnect_0_botao_s1_write_ports_inv <= not mm_interconnect_0_botao_s1_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_timestamp_timer_s1_write_ports_inv <= not mm_interconnect_0_timestamp_timer_s1_write;

	mm_interconnect_0_timer_geral_s1_write_ports_inv <= not mm_interconnect_0_timer_geral_s1_write;

	mm_interconnect_0_watchdog_timer_s1_write_ports_inv <= not mm_interconnect_0_watchdog_timer_s1_write;

	mm_interconnect_0_hex_0_s1_write_ports_inv <= not mm_interconnect_0_hex_0_s1_write;

	mm_interconnect_0_hex_5_s1_write_ports_inv <= not mm_interconnect_0_hex_5_s1_write;

	mm_interconnect_0_hex_4_s1_write_ports_inv <= not mm_interconnect_0_hex_4_s1_write;

	mm_interconnect_0_hex_3_s1_write_ports_inv <= not mm_interconnect_0_hex_3_s1_write;

	mm_interconnect_0_hex_2_s1_write_ports_inv <= not mm_interconnect_0_hex_2_s1_write;

	mm_interconnect_0_hex_1_s1_write_ports_inv <= not mm_interconnect_0_hex_1_s1_write;

	mm_interconnect_0_motor1_s1_write_ports_inv <= not mm_interconnect_0_motor1_s1_write;

	mm_interconnect_0_motor2_s1_write_ports_inv <= not mm_interconnect_0_motor2_s1_write;

	mm_interconnect_0_motor4_s1_write_ports_inv <= not mm_interconnect_0_motor4_s1_write;

	mm_interconnect_0_motor3_s1_write_ports_inv <= not mm_interconnect_0_motor3_s1_write;

	mm_interconnect_0_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_spi_control_port_read;

	mm_interconnect_0_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of sopc_2
