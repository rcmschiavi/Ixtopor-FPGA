// sopc_2.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module sopc_2 (
		input  wire [4:0] botoes_export,    //    botoes.export
		input  wire       clk_clk,          //       clk.clk
		input  wire [7:0] entrada_c_export, // entrada_c.export
		inout  wire [7:0] porta_a_export,   //   porta_a.export
		inout  wire [7:0] porta_b_export,   //   porta_b.export
		input  wire       reset_reset_n,    //     reset.reset_n
		output wire [7:0] saida_c_export,   //   saida_c.export
		input  wire       spi_MISO,         //       spi.MISO
		output wire       spi_MOSI,         //          .MOSI
		output wire       spi_SCLK,         //          .SCLK
		output wire [1:0] spi_SS_n,         //          .SS_n
		output wire       to_export,        //        to.export
		input  wire       uart_rxd,         //      uart.rxd
		output wire       uart_txd          //          .txd
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [17:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [17:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] mm_interconnect_0_adc_0_adc_slave_readdata;                // adc_0:readdata -> mm_interconnect_0:adc_0_adc_slave_readdata
	wire         mm_interconnect_0_adc_0_adc_slave_waitrequest;             // adc_0:waitrequest -> mm_interconnect_0:adc_0_adc_slave_waitrequest
	wire   [2:0] mm_interconnect_0_adc_0_adc_slave_address;                 // mm_interconnect_0:adc_0_adc_slave_address -> adc_0:address
	wire         mm_interconnect_0_adc_0_adc_slave_read;                    // mm_interconnect_0:adc_0_adc_slave_read -> adc_0:read
	wire         mm_interconnect_0_adc_0_adc_slave_write;                   // mm_interconnect_0:adc_0_adc_slave_write -> adc_0:write
	wire  [31:0] mm_interconnect_0_adc_0_adc_slave_writedata;               // mm_interconnect_0:adc_0_adc_slave_writedata -> adc_0:writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_memoria_s1_chipselect;                   // mm_interconnect_0:memoria_s1_chipselect -> memoria:chipselect
	wire  [31:0] mm_interconnect_0_memoria_s1_readdata;                     // memoria:readdata -> mm_interconnect_0:memoria_s1_readdata
	wire  [13:0] mm_interconnect_0_memoria_s1_address;                      // mm_interconnect_0:memoria_s1_address -> memoria:address
	wire   [3:0] mm_interconnect_0_memoria_s1_byteenable;                   // mm_interconnect_0:memoria_s1_byteenable -> memoria:byteenable
	wire         mm_interconnect_0_memoria_s1_write;                        // mm_interconnect_0:memoria_s1_write -> memoria:write
	wire  [31:0] mm_interconnect_0_memoria_s1_writedata;                    // mm_interconnect_0:memoria_s1_writedata -> memoria:writedata
	wire         mm_interconnect_0_memoria_s1_clken;                        // mm_interconnect_0:memoria_s1_clken -> memoria:clken
	wire         mm_interconnect_0_porta_a_s1_chipselect;                   // mm_interconnect_0:PORTA_A_s1_chipselect -> PORTA_A:chipselect
	wire  [31:0] mm_interconnect_0_porta_a_s1_readdata;                     // PORTA_A:readdata -> mm_interconnect_0:PORTA_A_s1_readdata
	wire   [2:0] mm_interconnect_0_porta_a_s1_address;                      // mm_interconnect_0:PORTA_A_s1_address -> PORTA_A:address
	wire         mm_interconnect_0_porta_a_s1_write;                        // mm_interconnect_0:PORTA_A_s1_write -> PORTA_A:write_n
	wire  [31:0] mm_interconnect_0_porta_a_s1_writedata;                    // mm_interconnect_0:PORTA_A_s1_writedata -> PORTA_A:writedata
	wire         mm_interconnect_0_porta_b_s1_chipselect;                   // mm_interconnect_0:PORTA_B_s1_chipselect -> PORTA_B:chipselect
	wire  [31:0] mm_interconnect_0_porta_b_s1_readdata;                     // PORTA_B:readdata -> mm_interconnect_0:PORTA_B_s1_readdata
	wire   [2:0] mm_interconnect_0_porta_b_s1_address;                      // mm_interconnect_0:PORTA_B_s1_address -> PORTA_B:address
	wire         mm_interconnect_0_porta_b_s1_write;                        // mm_interconnect_0:PORTA_B_s1_write -> PORTA_B:write_n
	wire  [31:0] mm_interconnect_0_porta_b_s1_writedata;                    // mm_interconnect_0:PORTA_B_s1_writedata -> PORTA_B:writedata
	wire         mm_interconnect_0_saida_c_s1_chipselect;                   // mm_interconnect_0:saida_C_s1_chipselect -> saida_C:chipselect
	wire  [31:0] mm_interconnect_0_saida_c_s1_readdata;                     // saida_C:readdata -> mm_interconnect_0:saida_C_s1_readdata
	wire   [1:0] mm_interconnect_0_saida_c_s1_address;                      // mm_interconnect_0:saida_C_s1_address -> saida_C:address
	wire         mm_interconnect_0_saida_c_s1_write;                        // mm_interconnect_0:saida_C_s1_write -> saida_C:write_n
	wire  [31:0] mm_interconnect_0_saida_c_s1_writedata;                    // mm_interconnect_0:saida_C_s1_writedata -> saida_C:writedata
	wire  [31:0] mm_interconnect_0_entrada_c_s1_readdata;                   // entrada_C:readdata -> mm_interconnect_0:entrada_C_s1_readdata
	wire   [1:0] mm_interconnect_0_entrada_c_s1_address;                    // mm_interconnect_0:entrada_C_s1_address -> entrada_C:address
	wire         mm_interconnect_0_uart_s1_chipselect;                      // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                        // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                         // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                            // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                   // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                           // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                       // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_botoes_s1_chipselect;                    // mm_interconnect_0:botoes_s1_chipselect -> botoes:chipselect
	wire  [31:0] mm_interconnect_0_botoes_s1_readdata;                      // botoes:readdata -> mm_interconnect_0:botoes_s1_readdata
	wire   [1:0] mm_interconnect_0_botoes_s1_address;                       // mm_interconnect_0:botoes_s1_address -> botoes:address
	wire         mm_interconnect_0_botoes_s1_write;                         // mm_interconnect_0:botoes_s1_write -> botoes:write_n
	wire  [31:0] mm_interconnect_0_botoes_s1_writedata;                     // mm_interconnect_0:botoes_s1_writedata -> botoes:writedata
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;             // mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;               // sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                // mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                  // mm_interconnect_0:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;              // mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_0_timestamp_timer_s1_chipselect;           // mm_interconnect_0:timestamp_timer_s1_chipselect -> timestamp_timer:chipselect
	wire  [15:0] mm_interconnect_0_timestamp_timer_s1_readdata;             // timestamp_timer:readdata -> mm_interconnect_0:timestamp_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timestamp_timer_s1_address;              // mm_interconnect_0:timestamp_timer_s1_address -> timestamp_timer:address
	wire         mm_interconnect_0_timestamp_timer_s1_write;                // mm_interconnect_0:timestamp_timer_s1_write -> timestamp_timer:write_n
	wire  [15:0] mm_interconnect_0_timestamp_timer_s1_writedata;            // mm_interconnect_0:timestamp_timer_s1_writedata -> timestamp_timer:writedata
	wire         mm_interconnect_0_timer_geral_s1_chipselect;               // mm_interconnect_0:timer_geral_s1_chipselect -> timer_geral:chipselect
	wire  [15:0] mm_interconnect_0_timer_geral_s1_readdata;                 // timer_geral:readdata -> mm_interconnect_0:timer_geral_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_geral_s1_address;                  // mm_interconnect_0:timer_geral_s1_address -> timer_geral:address
	wire         mm_interconnect_0_timer_geral_s1_write;                    // mm_interconnect_0:timer_geral_s1_write -> timer_geral:write_n
	wire  [15:0] mm_interconnect_0_timer_geral_s1_writedata;                // mm_interconnect_0:timer_geral_s1_writedata -> timer_geral:writedata
	wire         mm_interconnect_0_watchdog_timer_s1_chipselect;            // mm_interconnect_0:watchdog_timer_s1_chipselect -> watchdog_timer:chipselect
	wire  [15:0] mm_interconnect_0_watchdog_timer_s1_readdata;              // watchdog_timer:readdata -> mm_interconnect_0:watchdog_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_watchdog_timer_s1_address;               // mm_interconnect_0:watchdog_timer_s1_address -> watchdog_timer:address
	wire         mm_interconnect_0_watchdog_timer_s1_write;                 // mm_interconnect_0:watchdog_timer_s1_write -> watchdog_timer:write_n
	wire  [15:0] mm_interconnect_0_watchdog_timer_s1_writedata;             // mm_interconnect_0:watchdog_timer_s1_writedata -> watchdog_timer:writedata
	wire         mm_interconnect_0_spi_spi_control_port_chipselect;         // mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_readdata;           // spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_spi_control_port_address;            // mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	wire         mm_interconnect_0_spi_spi_control_port_read;               // mm_interconnect_0:spi_spi_control_port_read -> spi:read_n
	wire         mm_interconnect_0_spi_spi_control_port_write;              // mm_interconnect_0:spi_spi_control_port_write -> spi:write_n
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_writedata;          // mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // PORTA_B:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // spi:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // botoes:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // sys_clk_timer:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                  // timestamp_timer:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                  // timer_geral:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                  // watchdog_timer:irq -> irq_mapper:receiver8_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [PORTA_A:reset_n, PORTA_B:reset_n, botoes:reset_n, entrada_C:reset_n, jtag_uart:rst_n, memoria:reset, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, saida_C:reset_n, spi:reset_n, sys_clk_timer:reset_n, sysid:reset_n, timer_geral:reset_n, timestamp_timer:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [memoria:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [adc_0:reset, mm_interconnect_0:adc_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset, watchdog_timer:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                    // rst_controller_002:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	wire         watchdog_timer_resetrequest_reset;                         // watchdog_timer:resetrequest -> rst_controller_002:reset_in2

	sopc_2_PORTA_A porta_a (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_porta_a_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_porta_a_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_porta_a_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_porta_a_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_porta_a_s1_readdata),   //                    .readdata
		.bidir_port (porta_a_export)                           // external_connection.export
	);

	sopc_2_PORTA_B porta_b (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_porta_b_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_porta_b_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_porta_b_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_porta_b_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_porta_b_s1_readdata),   //                    .readdata
		.bidir_port (porta_b_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	sopc_2_adc_0 #(
		.board          ("DE10-Lite"),
		.board_rev      ("Autodetect"),
		.tsclk          (5),
		.numch          (5),
		.max10pllmultby (1),
		.max10plldivby  (5)
	) adc_0 (
		.clock       (clk_clk),                                       //       clk.clk
		.reset       (rst_controller_001_reset_out_reset),            //     reset.reset
		.write       (mm_interconnect_0_adc_0_adc_slave_write),       // adc_slave.write
		.readdata    (mm_interconnect_0_adc_0_adc_slave_readdata),    //          .readdata
		.writedata   (mm_interconnect_0_adc_0_adc_slave_writedata),   //          .writedata
		.address     (mm_interconnect_0_adc_0_adc_slave_address),     //          .address
		.waitrequest (mm_interconnect_0_adc_0_adc_slave_waitrequest), //          .waitrequest
		.read        (mm_interconnect_0_adc_0_adc_slave_read),        //          .read
		.adc_sclk    (),                                              // (terminated)
		.adc_cs_n    (),                                              // (terminated)
		.adc_dout    (1'b0),                                          // (terminated)
		.adc_din     ()                                               // (terminated)
	);

	sopc_2_botoes botoes (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_botoes_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_botoes_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_botoes_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_botoes_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_botoes_s1_readdata),   //                    .readdata
		.in_port    (botoes_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                //                 irq.irq
	);

	sopc_2_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	sopc_2_entrada_C entrada_c (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_entrada_c_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_entrada_c_s1_readdata), //                    .readdata
		.in_port  (entrada_c_export)                         // external_connection.export
	);

	sopc_2_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	sopc_2_memoria memoria (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_memoria_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoria_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoria_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoria_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoria_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoria_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoria_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	sopc_2_saida_C saida_c (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_saida_c_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_saida_c_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_saida_c_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_saida_c_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_saida_c_s1_readdata),   //                    .readdata
		.out_port   (saida_c_export)                           // external_connection.export
	);

	sopc_2_spi spi (
		.clk           (clk_clk),                                           //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                          //              irq.irq
		.MISO          (spi_MISO),                                          //         external.export
		.MOSI          (spi_MOSI),                                          //                 .export
		.SCLK          (spi_SCLK),                                          //                 .export
		.SS_n          (spi_SS_n)                                           //                 .export
	);

	sopc_2_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                       //   irq.irq
	);

	sopc_2_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	sopc_2_timer_geral timer_geral (
		.clk           (clk_clk),                                     //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),             //         reset.reset_n
		.address       (mm_interconnect_0_timer_geral_s1_address),    //            s1.address
		.writedata     (mm_interconnect_0_timer_geral_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_0_timer_geral_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_0_timer_geral_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_0_timer_geral_s1_write),     //              .write_n
		.irq           (irq_mapper_receiver7_irq),                    //           irq.irq
		.timeout_pulse (to_export)                                    // external_port.export
	);

	sopc_2_timestamp_timer timestamp_timer (
		.clk        (clk_clk),                                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 // reset.reset_n
		.address    (mm_interconnect_0_timestamp_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                         //   irq.irq
	);

	sopc_2_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	sopc_2_watchdog_timer watchdog_timer (
		.clk          (clk_clk),                                        //          clk.clk
		.reset_n      (~rst_controller_002_reset_out_reset),            //        reset.reset_n
		.address      (mm_interconnect_0_watchdog_timer_s1_address),    //           s1.address
		.writedata    (mm_interconnect_0_watchdog_timer_s1_writedata),  //             .writedata
		.readdata     (mm_interconnect_0_watchdog_timer_s1_readdata),   //             .readdata
		.chipselect   (mm_interconnect_0_watchdog_timer_s1_chipselect), //             .chipselect
		.write_n      (~mm_interconnect_0_watchdog_timer_s1_write),     //             .write_n
		.irq          (irq_mapper_receiver8_irq),                       //          irq.irq
		.resetrequest (watchdog_timer_resetrequest_reset)               // resetrequest.reset
	);

	sopc_2_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                 (clk_clk),                                                   //                               clk_clk.clk
		.adc_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                        //     adc_0_reset_reset_bridge_in_reset.reset
		.cpu_reset_reset_bridge_in_reset_reset       (rst_controller_002_reset_out_reset),                        //       cpu_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // jtag_uart_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                     (cpu_data_master_address),                                   //                       cpu_data_master.address
		.cpu_data_master_waitrequest                 (cpu_data_master_waitrequest),                               //                                      .waitrequest
		.cpu_data_master_byteenable                  (cpu_data_master_byteenable),                                //                                      .byteenable
		.cpu_data_master_read                        (cpu_data_master_read),                                      //                                      .read
		.cpu_data_master_readdata                    (cpu_data_master_readdata),                                  //                                      .readdata
		.cpu_data_master_write                       (cpu_data_master_write),                                     //                                      .write
		.cpu_data_master_writedata                   (cpu_data_master_writedata),                                 //                                      .writedata
		.cpu_data_master_debugaccess                 (cpu_data_master_debugaccess),                               //                                      .debugaccess
		.cpu_instruction_master_address              (cpu_instruction_master_address),                            //                cpu_instruction_master.address
		.cpu_instruction_master_waitrequest          (cpu_instruction_master_waitrequest),                        //                                      .waitrequest
		.cpu_instruction_master_read                 (cpu_instruction_master_read),                               //                                      .read
		.cpu_instruction_master_readdata             (cpu_instruction_master_readdata),                           //                                      .readdata
		.adc_0_adc_slave_address                     (mm_interconnect_0_adc_0_adc_slave_address),                 //                       adc_0_adc_slave.address
		.adc_0_adc_slave_write                       (mm_interconnect_0_adc_0_adc_slave_write),                   //                                      .write
		.adc_0_adc_slave_read                        (mm_interconnect_0_adc_0_adc_slave_read),                    //                                      .read
		.adc_0_adc_slave_readdata                    (mm_interconnect_0_adc_0_adc_slave_readdata),                //                                      .readdata
		.adc_0_adc_slave_writedata                   (mm_interconnect_0_adc_0_adc_slave_writedata),               //                                      .writedata
		.adc_0_adc_slave_waitrequest                 (mm_interconnect_0_adc_0_adc_slave_waitrequest),             //                                      .waitrequest
		.botoes_s1_address                           (mm_interconnect_0_botoes_s1_address),                       //                             botoes_s1.address
		.botoes_s1_write                             (mm_interconnect_0_botoes_s1_write),                         //                                      .write
		.botoes_s1_readdata                          (mm_interconnect_0_botoes_s1_readdata),                      //                                      .readdata
		.botoes_s1_writedata                         (mm_interconnect_0_botoes_s1_writedata),                     //                                      .writedata
		.botoes_s1_chipselect                        (mm_interconnect_0_botoes_s1_chipselect),                    //                                      .chipselect
		.cpu_debug_mem_slave_address                 (mm_interconnect_0_cpu_debug_mem_slave_address),             //                   cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                   (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                      .write
		.cpu_debug_mem_slave_read                    (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                      .read
		.cpu_debug_mem_slave_readdata                (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                      .readdata
		.cpu_debug_mem_slave_writedata               (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                      .writedata
		.cpu_debug_mem_slave_byteenable              (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                      .byteenable
		.cpu_debug_mem_slave_waitrequest             (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                      .waitrequest
		.cpu_debug_mem_slave_debugaccess             (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                      .debugaccess
		.entrada_C_s1_address                        (mm_interconnect_0_entrada_c_s1_address),                    //                          entrada_C_s1.address
		.entrada_C_s1_readdata                       (mm_interconnect_0_entrada_c_s1_readdata),                   //                                      .readdata
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.memoria_s1_address                          (mm_interconnect_0_memoria_s1_address),                      //                            memoria_s1.address
		.memoria_s1_write                            (mm_interconnect_0_memoria_s1_write),                        //                                      .write
		.memoria_s1_readdata                         (mm_interconnect_0_memoria_s1_readdata),                     //                                      .readdata
		.memoria_s1_writedata                        (mm_interconnect_0_memoria_s1_writedata),                    //                                      .writedata
		.memoria_s1_byteenable                       (mm_interconnect_0_memoria_s1_byteenable),                   //                                      .byteenable
		.memoria_s1_chipselect                       (mm_interconnect_0_memoria_s1_chipselect),                   //                                      .chipselect
		.memoria_s1_clken                            (mm_interconnect_0_memoria_s1_clken),                        //                                      .clken
		.PORTA_A_s1_address                          (mm_interconnect_0_porta_a_s1_address),                      //                            PORTA_A_s1.address
		.PORTA_A_s1_write                            (mm_interconnect_0_porta_a_s1_write),                        //                                      .write
		.PORTA_A_s1_readdata                         (mm_interconnect_0_porta_a_s1_readdata),                     //                                      .readdata
		.PORTA_A_s1_writedata                        (mm_interconnect_0_porta_a_s1_writedata),                    //                                      .writedata
		.PORTA_A_s1_chipselect                       (mm_interconnect_0_porta_a_s1_chipselect),                   //                                      .chipselect
		.PORTA_B_s1_address                          (mm_interconnect_0_porta_b_s1_address),                      //                            PORTA_B_s1.address
		.PORTA_B_s1_write                            (mm_interconnect_0_porta_b_s1_write),                        //                                      .write
		.PORTA_B_s1_readdata                         (mm_interconnect_0_porta_b_s1_readdata),                     //                                      .readdata
		.PORTA_B_s1_writedata                        (mm_interconnect_0_porta_b_s1_writedata),                    //                                      .writedata
		.PORTA_B_s1_chipselect                       (mm_interconnect_0_porta_b_s1_chipselect),                   //                                      .chipselect
		.saida_C_s1_address                          (mm_interconnect_0_saida_c_s1_address),                      //                            saida_C_s1.address
		.saida_C_s1_write                            (mm_interconnect_0_saida_c_s1_write),                        //                                      .write
		.saida_C_s1_readdata                         (mm_interconnect_0_saida_c_s1_readdata),                     //                                      .readdata
		.saida_C_s1_writedata                        (mm_interconnect_0_saida_c_s1_writedata),                    //                                      .writedata
		.saida_C_s1_chipselect                       (mm_interconnect_0_saida_c_s1_chipselect),                   //                                      .chipselect
		.spi_spi_control_port_address                (mm_interconnect_0_spi_spi_control_port_address),            //                  spi_spi_control_port.address
		.spi_spi_control_port_write                  (mm_interconnect_0_spi_spi_control_port_write),              //                                      .write
		.spi_spi_control_port_read                   (mm_interconnect_0_spi_spi_control_port_read),               //                                      .read
		.spi_spi_control_port_readdata               (mm_interconnect_0_spi_spi_control_port_readdata),           //                                      .readdata
		.spi_spi_control_port_writedata              (mm_interconnect_0_spi_spi_control_port_writedata),          //                                      .writedata
		.spi_spi_control_port_chipselect             (mm_interconnect_0_spi_spi_control_port_chipselect),         //                                      .chipselect
		.sys_clk_timer_s1_address                    (mm_interconnect_0_sys_clk_timer_s1_address),                //                      sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                      (mm_interconnect_0_sys_clk_timer_s1_write),                  //                                      .write
		.sys_clk_timer_s1_readdata                   (mm_interconnect_0_sys_clk_timer_s1_readdata),               //                                      .readdata
		.sys_clk_timer_s1_writedata                  (mm_interconnect_0_sys_clk_timer_s1_writedata),              //                                      .writedata
		.sys_clk_timer_s1_chipselect                 (mm_interconnect_0_sys_clk_timer_s1_chipselect),             //                                      .chipselect
		.sysid_control_slave_address                 (mm_interconnect_0_sysid_control_slave_address),             //                   sysid_control_slave.address
		.sysid_control_slave_readdata                (mm_interconnect_0_sysid_control_slave_readdata),            //                                      .readdata
		.timer_geral_s1_address                      (mm_interconnect_0_timer_geral_s1_address),                  //                        timer_geral_s1.address
		.timer_geral_s1_write                        (mm_interconnect_0_timer_geral_s1_write),                    //                                      .write
		.timer_geral_s1_readdata                     (mm_interconnect_0_timer_geral_s1_readdata),                 //                                      .readdata
		.timer_geral_s1_writedata                    (mm_interconnect_0_timer_geral_s1_writedata),                //                                      .writedata
		.timer_geral_s1_chipselect                   (mm_interconnect_0_timer_geral_s1_chipselect),               //                                      .chipselect
		.timestamp_timer_s1_address                  (mm_interconnect_0_timestamp_timer_s1_address),              //                    timestamp_timer_s1.address
		.timestamp_timer_s1_write                    (mm_interconnect_0_timestamp_timer_s1_write),                //                                      .write
		.timestamp_timer_s1_readdata                 (mm_interconnect_0_timestamp_timer_s1_readdata),             //                                      .readdata
		.timestamp_timer_s1_writedata                (mm_interconnect_0_timestamp_timer_s1_writedata),            //                                      .writedata
		.timestamp_timer_s1_chipselect               (mm_interconnect_0_timestamp_timer_s1_chipselect),           //                                      .chipselect
		.uart_s1_address                             (mm_interconnect_0_uart_s1_address),                         //                               uart_s1.address
		.uart_s1_write                               (mm_interconnect_0_uart_s1_write),                           //                                      .write
		.uart_s1_read                                (mm_interconnect_0_uart_s1_read),                            //                                      .read
		.uart_s1_readdata                            (mm_interconnect_0_uart_s1_readdata),                        //                                      .readdata
		.uart_s1_writedata                           (mm_interconnect_0_uart_s1_writedata),                       //                                      .writedata
		.uart_s1_begintransfer                       (mm_interconnect_0_uart_s1_begintransfer),                   //                                      .begintransfer
		.uart_s1_chipselect                          (mm_interconnect_0_uart_s1_chipselect),                      //                                      .chipselect
		.watchdog_timer_s1_address                   (mm_interconnect_0_watchdog_timer_s1_address),               //                     watchdog_timer_s1.address
		.watchdog_timer_s1_write                     (mm_interconnect_0_watchdog_timer_s1_write),                 //                                      .write
		.watchdog_timer_s1_readdata                  (mm_interconnect_0_watchdog_timer_s1_readdata),              //                                      .readdata
		.watchdog_timer_s1_writedata                 (mm_interconnect_0_watchdog_timer_s1_writedata),             //                                      .writedata
		.watchdog_timer_s1_chipselect                (mm_interconnect_0_watchdog_timer_s1_chipselect)             //                                      .chipselect
	);

	sopc_2_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),           // receiver8.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.reset_in2      (watchdog_timer_resetrequest_reset),      // reset_in2.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
